module bus_top (

);

endmodule
