library verilog;
use verilog.vl_types.all;
entity ex is
    port(
        rst             : in     vl_logic;
        aluop_i         : in     vl_logic_vector(7 downto 0);
        alusel_i        : in     vl_logic_vector(2 downto 0);
        reg1_i          : in     vl_logic_vector(31 downto 0);
        reg2_i          : in     vl_logic_vector(31 downto 0);
        wd_i            : in     vl_logic_vector(4 downto 0);
        wreg_i          : in     vl_logic;
        inst_i          : in     vl_logic_vector(31 downto 0);
        excepttype_i    : in     vl_logic_vector(31 downto 0);
        current_inst_address_i: in     vl_logic_vector(31 downto 0);
        hi_i            : in     vl_logic_vector(31 downto 0);
        lo_i            : in     vl_logic_vector(31 downto 0);
        wb_hi_i         : in     vl_logic_vector(31 downto 0);
        wb_lo_i         : in     vl_logic_vector(31 downto 0);
        wb_whilo_i      : in     vl_logic;
        mem_hi_i        : in     vl_logic_vector(31 downto 0);
        mem_lo_i        : in     vl_logic_vector(31 downto 0);
        mem_whilo_i     : in     vl_logic;
        hilo_temp_i     : in     vl_logic_vector(63 downto 0);
        cnt_i           : in     vl_logic_vector(1 downto 0);
        link_address_i  : in     vl_logic_vector(31 downto 0);
        is_in_delayslot_i: in     vl_logic;
        mem_cp0_reg_we  : in     vl_logic;
        mem_cp0_reg_write_addr: in     vl_logic_vector(4 downto 0);
        mem_cp0_reg_data: in     vl_logic_vector(31 downto 0);
        wb_cp0_reg_we   : in     vl_logic;
        wb_cp0_reg_write_addr: in     vl_logic_vector(4 downto 0);
        wb_cp0_reg_data : in     vl_logic_vector(31 downto 0);
        cp0_reg_data_i  : in     vl_logic_vector(31 downto 0);
        cp0_reg_read_addr_o: out    vl_logic_vector(4 downto 0);
        cp0_reg_we_o    : out    vl_logic;
        cp0_reg_write_addr_o: out    vl_logic_vector(4 downto 0);
        cp0_reg_data_o  : out    vl_logic_vector(31 downto 0);
        wd_o            : out    vl_logic_vector(4 downto 0);
        wreg_o          : out    vl_logic;
        wdata_o         : out    vl_logic_vector(31 downto 0);
        hi_o            : out    vl_logic_vector(31 downto 0);
        lo_o            : out    vl_logic_vector(31 downto 0);
        whilo_o         : out    vl_logic;
        hilo_temp_o     : out    vl_logic_vector(63 downto 0);
        cnt_o           : out    vl_logic_vector(1 downto 0);
        excepttype_o    : out    vl_logic_vector(31 downto 0);
        is_in_delayslot_o: out    vl_logic;
        current_inst_address_o: out    vl_logic_vector(31 downto 0);
        aluop_o         : out    vl_logic_vector(7 downto 0);
        mem_addr_o      : out    vl_logic_vector(31 downto 0);
        reg2_o          : out    vl_logic_vector(31 downto 0);
        stallreq        : out    vl_logic
    );
end ex;
