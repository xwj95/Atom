module ram (
	input bus_clk_i,
	input bus_rst_i,
	input [31:0] bus_addr_i,
	input [31:0] bus_data_i,
	output reg[31:0] bus_data_o,
	input bus_select_i,
	input bus_we_i,
	output bus_ack_o,

	output [19:0] baseram_addr,
	inout [31:0] baseram_data,
	output baseram_ce,
	output baseram_oe,
	output baseram_we,

	output [19:0] extram_addr,
	inout [31:0] extram_data,
	output extram_ce,
	output extram_oe,
	output extram_we
	);

	ram_driver ram_driver_inst (
		bus_clk_i, bus_rst_i, 
		bus_select_i, !bus_we_i, bus_we_i, 
		{bus_addr_i[19], bus_addr_i[19:0]}, bus_data_i, bus_data_o,
		baseram_addr, baseram_data, 
		baseram_ce, baseram_oe, baseram_we, 
		extram_addr, extram_data, 
		extram_ce, extram_oe, extram_we, bus_ack_o
	);

endmodule
