`include "defines.v"

module wishbone_bus(
	input		wire					clk,
	input		wire					rst,

	//来自ctrl模块
	input		wire[5:0]				stall_i,
	input		wire					flush_i,

	//CPU侧的接口
	input		wire					cpu_ce_i,
	input		wire[`RegBus]			cpu_data_i,
	input		wire[`RegBus]			cpu_addr_i,
	input		wire					cpu_we_i,
	input		wire[3:0]				cpu_sel_i,
	output		reg[`RegBus]			cpu_data_o,

	//Wishbone侧的接口
	input		wire[`RegBus]			wishbone_data_i,
	input		wire					wishbone_ack_i,
	output		reg[`RegBus]			wishbone_addr_o,
	output		reg[`RegBus]			wishbone_data_o,
	output		reg						wishbone_we_o,
	output		reg[3:0]				wishbone_sel_o,
	output		reg						wishbone_stb_o,
	output		reg						wishbone_cyc_o,

	output		reg						stallreq
	);

	reg[1:0] wishbone_state;			//保存Wishbone总线接口模块的状态
	reg[`RegBus] rd_buf;				//寄存通过Wishbone总线访问到的数据

	/*********************		第一段：控制状态转化的时序电路		*********************/
	always @ (posedge clk) begin
		if (rst == `RstEnable) begin
			wishbone_state <= `WB_IDLE;
			wishbone_addr_o <= `ZeroWord;
			wishbone_data_o <= `ZeroWord;
			wishbone_we_o <= `WriteDisable;
			wishbone_sel_o <= 4'b0000;
			wishbone_stb_o <= 1'b0;
			wishbone_cyc_o <= 1'b0;
			rd_buf <= `ZeroWord;
		end else begin
			case (wishbone_state)
				`WB_IDLE: begin								//WB_IDLE状态
					if ((cpu_ce_i == 1'b1) && (flush_i == `False_v)) begin
						wishbone_stb_o <= 1'b1;
						wishbone_cyc_o <= 1'b1;
						wishbone_addr_o <= cpu_addr_i;
						wishbone_data_o <= cpu_data_i;
						wishbone_we_o <= cpu_we_i;
						wishbone_sel_o <= cpu_sel_i;
						wishbone_state <= `WB_BUSY;			//进入WB_BUSY状态
					end
				end
				`WB_BUSY: begin								//WB_BUSY状态
					if (wishbone_ack_i == 1'b1) begin
						wishbone_stb_o <= 1'b0;
						wishbone_cyc_o <= 1'b0;
						wishbone_addr_o <= `ZeroWord;
						wishbone_data_o <= `ZeroWord;
						wishbone_we_o <= `WriteDisable;
						wishbone_sel_o <= 4'b0000;
						wishbone_state <= `WB_IDLE;
						if (cpu_we_i == `WriteDisable) begin
							rd_buf <= wishbone_data_i;
						end
						if (stall_i != 6'b000000) begin		//进入WB_WAIT_FOR_STALL状态
							wishbone_state <= `WB_WAIT_FOR_STALL;
						end
					end else if (flush_i == `True_v) begin
						wishbone_stb_o <= 1'b0;
						wishbone_cyc_o <= 1'b0;
						wishbone_addr_o <= `ZeroWord;
						wishbone_data_o <= `ZeroWord;
						wishbone_we_o <= `WriteDisable;
						wishbone_sel_o <= 4'b0000;
						wishbone_state <= `WB_IDLE;			//进入WB_IDLE状态
						rd_buf <= `ZeroWord;
					end
				end
				`WB_WAIT_FOR_STALL: begin					//WB_WAIT_FOR_STALL状态
					if (stall_i == 6'b000000) begin
						wishbone_state <= `WB_IDLE;			//进入WB_IDLE状态
					end
				end
				default: begin
				end
			endcase
		end
	end

	/*********************		第二段：给处理器接口信号赋值的组合电路		*********************/
	always @ (*) begin
		if (rst == `RstEnable) begin
			stallreq <= `NoStop;
			cpu_data_o <= `ZeroWord;
		end else begin
			stallreq <= `NoStop;
			case (wishbone_state)
				`WB_IDLE: begin								//WB_IDLE状态
					if ((cpu_ce_i == 1'b1) && (flush_i == `False_v)) begin
						stallreq <= `Stop;
						cpu_data_o <= `ZeroWord;
					end
				end
				`WB_BUSY: begin								//WB_BUSY状态
					if (wishbone_ack_i == 1'b1) begin
						stallreq <= `NoStop;
						if (wishbone_we_o == `WriteDisable) begin
							cpu_data_o <= wishbone_data_i;
						end else begin
							cpu_data_o <= `ZeroWord;
						end
					end else begin
						stallreq <= `Stop;
						cpu_data_o <= `ZeroWord;
					end
				end
				`WB_WAIT_FOR_STALL: begin					//WB_WAIT_FOR_STALL状态
					stallreq <= `NoStop;
					cpu_data_o <= rd_buf;
				end
				default: begin
				end
			endcase
		end
	end

endmodule
