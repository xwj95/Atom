library verilog;
use verilog.vl_types.all;
entity ASSERTION_ERROR is
    port(
        param           : in     vl_logic
    );
end ASSERTION_ERROR;
